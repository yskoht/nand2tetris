localparam H_PERIOD = 10'd800;
localparam H_FRONT = 10'd16;
localparam H_WIDTH = 10'd96;
localparam H_BACK = 10'd48;

localparam V_PERIOD = 10'd525;
localparam V_FRONT = 10'd10;
localparam V_WIDTH = 10'd2;
localparam V_BACK = 10'd33;
